import cds_rnm_pkg::*;

package nettypes_pkg;

  nettype wreal1driver voltage_net;

endpackage
